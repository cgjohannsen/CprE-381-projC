libray IEEE;
use IEEE.std_logic_1164.all

entity IF_ID is 
    port ();

end IF_ID;

architecture struct of IF_ID is

end struct;